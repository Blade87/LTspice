.SUBCKT C0402C104K3PAC 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 10000 Hz
*KEMET Model RLC Cerm
R1 3 4 3.78656268119812
R2 2 5 1.50999999046326
R3 1 6 11109999616
L1 1 2 1.19999996051057E-11
L2 2 3 2.27999992497008E-10
C1 4 6 8.73000018941639E-08
C2 5 6 3.90000009536743E-12
.ENDS